`ifdef VERILATE
    localparam FILE_PATH = "D:/sysI/sys1-sp25/repo/sys-project/lab3-3/syn/initial.hex";
`else
    localparam FILE_PATH = "D:/sysI/sys1-sp25/repo/sys-project/lab3-3/syn/initial.hex";
`endif